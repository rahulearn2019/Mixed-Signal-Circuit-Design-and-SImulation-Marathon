* /home/tiw.rahul45/eSim-2.3/library/SubcircuitLibrary/rahul_inv/rahul_inv.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Fri 07 Oct 2022 11:13:02 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v1  Net-_SC1-Pad3_ GND DC		
SC2  Net-_SC1-Pad1_ Net-_SC1-Pad2_ GND GND sky130_fd_pr__nfet_01v8		
SC1  Net-_SC1-Pad1_ Net-_SC1-Pad2_ Net-_SC1-Pad3_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8		
U2  Net-_SC1-Pad2_ Net-_SC1-Pad1_ PORT		

.end
